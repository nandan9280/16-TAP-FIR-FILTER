module ripple_carry_adder_32bit(A, B, Cin, Sum);
    input [31:0] A, B;
    input Cin;
    output [31:0] Sum;
    wire [31:0] carry;

    full_adder FA0(A[0], B[0], Cin, Sum[0], carry[0]);
    full_adder FA1(A[1], B[1], carry[0], Sum[1], carry[1]);
    full_adder FA2(A[2], B[2], carry[1], Sum[2], carry[2]);
    full_adder FA3(A[3], B[3], carry[2], Sum[3], carry[3]);
    full_adder FA4(A[4], B[4], carry[3], Sum[4], carry[4]);
    full_adder FA5(A[5], B[5], carry[4], Sum[5], carry[5]);
    full_adder FA6(A[6], B[6], carry[5], Sum[6], carry[6]);
    full_adder FA7(A[7], B[7], carry[6], Sum[7], carry[7]);
    full_adder FA8(A[8], B[8], carry[7], Sum[8], carry[8]);
    full_adder FA9(A[9], B[9], carry[8], Sum[9], carry[9]);
    full_adder FA10(A[10], B[10], carry[9], Sum[10], carry[10]);
    full_adder FA11(A[11], B[11], carry[10], Sum[11], carry[11]);
    full_adder FA12(A[12], B[12], carry[11], Sum[12], carry[12]);
    full_adder FA13(A[13], B[13], carry[12], Sum[13], carry[13]);
    full_adder FA14(A[14], B[14], carry[13], Sum[14], carry[14]);
    full_adder FA15(A[15], B[15], carry[14], Sum[15], carry[15]);
    full_adder FA16(A[16], B[16], carry[15], Sum[16], carry[16]);
    full_adder FA17(A[17], B[17], carry[16], Sum[17], carry[17]);
    full_adder FA18(A[18], B[18], carry[17], Sum[18], carry[18]);
    full_adder FA19(A[19], B[19], carry[18], Sum[19], carry[19]);
    full_adder FA20(A[20], B[20], carry[19], Sum[20], carry[20]);
    full_adder FA21(A[21], B[21], carry[20], Sum[21], carry[21]);
    full_adder FA22(A[22], B[22], carry[21], Sum[22], carry[22]);
    full_adder FA23(A[23], B[23], carry[22], Sum[23], carry[23]);
    full_adder FA24(A[24], B[24], carry[23], Sum[24], carry[24]);
    full_adder FA25(A[25], B[25], carry[24], Sum[25], carry[25]);
    full_adder FA26(A[26], B[26], carry[25], Sum[26], carry[26]);
    full_adder FA27(A[27], B[27], carry[26], Sum[27], carry[27]);
    full_adder FA28(A[28], B[28], carry[27], Sum[28], carry[28]);
    full_adder FA29(A[29], B[29], carry[28], Sum[29], carry[29]);
    full_adder FA30(A[30], B[30], carry[29], Sum[30], carry[30]);
    full_adder FA31(A[31], B[31], carry[30], Sum[31], carry[31]);
endmodule